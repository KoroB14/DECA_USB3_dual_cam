//////////////////////////////////////////////////////////////////////////////////
// Dmitry Koroteev
// korob14@gmail.com
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module MainFSM
#(	//Image params
	parameter IM_X = 1280,
	parameter IM_Y = 720,
	parameter COLOR_MODE = 2
)

(
    input 					USB_CLK,
	 input 					rst_n,
    input 					DMA0_Ready,
	 input 					DMA0_Watermark,
	 input 					DMA1_Ready, 
	 input 					DMA1_Watermark, 
	 output reg 			WR, 
	 output reg 			RD,
	 output reg 			LastWRData,
	 output reg 			OE,
	 output reg	[1:0]		DMA0_Address,
	 inout 		[15:0] 	DQ,
	 
	 //Cam interfaces
	 Cam_If.Cons 			Cam_R_IF,
	 Cam_If.Cons 			Cam_L_IF
);



//FIFO params
localparam BYTE_MUL = 'd2;
localparam BYTES = COLOR_MODE * IM_X + 2;
localparam WORDS = BYTES / BYTE_MUL;
localparam XWORDS = $clog2(2*WORDS);
//Packet params
localparam PacketID = (COLOR_MODE == 1) ? 16'h01AA : ((COLOR_MODE == 2) ? 16'h01BB : 0);
//Ctrl params
localparam GET_CFG = 8'h01;
localparam STRT_ST = 8'h11;
localparam STOP_ST = 8'h0f;

//FSM states
enum logic [10:0] {	WAIT4DMA 	= 11'b00000000001,
							WRITE,
							PAUSE_W,
							DR_READ,
							READ,
							PAUSE_R,
							RD_CMD,
							SEND_CFG,
							START_ST,
							STP_ST,
							SW_BUF} CurrentState, NextState;

//declarations
reg DMA0_Ready_t, DMA0_Watermark_t, DMA0_Ready_r, DMA0_Watermark_r, DMA1_Ready_r, DMA1_Watermark_r;							
reg [15:0] DATA_IN, DATA;
reg [15:0] pkt_data;
reg [2:0] lat_count;
reg [15:0] send_cnt;
reg [15:0] line_cnt_r, line_cnt_l;
reg [1:0] rdaddress;
reg start_stream;
wire rdreq_r, rdreq_l, rdreq;
wire [15:0] fifo_data_r, fifo_data_l;
wire fifo_full_r, fifo_full_l;
wire fifo_empty_r, fifo_empty_l;
wire [XWORDS - 1 : 0] usedw_r, usedw_l, usedw, usedw_other;
wire start_cond;
//assignments
assign DQ = WR ? DATA : 16'hzzzz;
assign Cam_R_IF.out_ready = ~fifo_full_r;
assign Cam_L_IF.out_ready = ~fifo_full_l;
assign Cam_R_IF.start_stream = start_stream;
assign Cam_L_IF.start_stream = start_stream;

//reg DMA flags
always @ (posedge USB_CLK)
begin
	{DMA0_Ready_t, DMA0_Watermark_t, DMA1_Ready_r, DMA1_Watermark_r} <= {DMA0_Ready, DMA0_Watermark, DMA1_Ready, DMA1_Watermark};
	{DMA0_Ready_r, DMA0_Watermark_r} <= {DMA0_Ready_t, DMA0_Watermark_t};
end

//reg input data
always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n) 	
	DATA_IN <= 0;
else 
	if (CurrentState == READ) 
		DATA_IN <= DQ;

//FIFO Right
dc_data_fifo 
#(.ADDR_W(XWORDS),
  .DATA_IN_W(8),
  .DATA_OUT_W(8*BYTE_MUL)) 
dc_data_fifo_r
(
	.rdclk(USB_CLK),
	.wrclk(Cam_R_IF.PCLK_cam),
	.rst_n(rst_n & start_stream),
	.rdreq(rdreq_r & !fifo_empty_r),
	.wrreq(Cam_R_IF.pixel_valid & !fifo_full_r),
	.data_in(Cam_R_IF.pixel),
	.data_out(fifo_data_r),
	.rdempty(fifo_empty_r),
	.wrfull(fifo_full_r),
	.rdusedw(usedw_r)
);

//FIFO Left
dc_data_fifo 
#(.ADDR_W(XWORDS),
  .DATA_IN_W(8),
  .DATA_OUT_W(8*BYTE_MUL)) 
dc_data_fifo_l
(
	.rdclk(USB_CLK),
	.wrclk(Cam_L_IF.PCLK_cam),
	.rst_n(rst_n & start_stream),
	.rdreq(rdreq_l & !fifo_empty_l),
	.wrreq(Cam_L_IF.pixel_valid & !fifo_full_l),
	.data_in(Cam_L_IF.pixel),
	.data_out(fifo_data_l),
	.rdempty(fifo_empty_l),
	.wrfull(fifo_full_l),
	.rdusedw(usedw_l)
);

//Stream params rom
always @(*)
case(rdaddress)
	'h00	:	pkt_data = PacketID; // Packet ID
	'h01	: 	pkt_data = IM_X; // IM_X
	'h02	: 	pkt_data = IM_Y; // IM_Y
	default: pkt_data = 8'h00;
endcase

always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n)
	rdaddress <= 0;
else if (CurrentState == SEND_CFG)
	rdaddress <= rdaddress + 1'b1;
else
	rdaddress <= 0;

//Control signals
always @ (posedge USB_CLK) 
begin
	 WR <= (CurrentState == WRITE) || (CurrentState == SEND_CFG) ;
	 LastWRData <= (rdaddress == 'h02) && (CurrentState == SEND_CFG);
	 RD <= (CurrentState == DR_READ) && (lat_count == 1);
	 OE <= (CurrentState == DR_READ) || (CurrentState == READ);
	 DMA0_Address[1] <= (CurrentState == DR_READ) || (CurrentState == READ);
end

//Data mux
always @ (posedge USB_CLK) 
if (((CurrentState == WRITE) || (CurrentState == PAUSE_W)) && (send_cnt == 0))
		DATA <= DMA0_Address[0] ? line_cnt_l : line_cnt_r;
else if (CurrentState == SEND_CFG)
		DATA <= pkt_data;
else
		DATA <= DMA0_Address[0] ? fifo_data_l : fifo_data_r;


//reg start_stream;
always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n)
	start_stream <= 0;
else if (CurrentState == START_ST)
	start_stream <= 1'b1;
else if (CurrentState == STP_ST)
	start_stream <= 0;

//FSM state
always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n) 
	CurrentState <= WAIT4DMA;
else 
	CurrentState <= NextState;

//latency counter
always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n)
	lat_count <= 0;
else if ((CurrentState == DR_READ) || (CurrentState == PAUSE_R) || (CurrentState == PAUSE_W) || (CurrentState == SW_BUF))
	lat_count <= lat_count + 1'b1;
else 
	lat_count <= 0;
	
//fifo selector
always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n)
	DMA0_Address[0] <= 0;
else if ((CurrentState == SW_BUF) && (lat_count == 0))
	DMA0_Address[0] <= ~DMA0_Address[0];

assign rdreq = (CurrentState == WRITE) && ((send_cnt <= WORDS - 2));
assign rdreq_r = rdreq  && !DMA0_Address[0]; 
assign rdreq_l = rdreq && DMA0_Address[0];
assign usedw = DMA0_Address[0] ? usedw_l : usedw_r;	
assign usedw_other = DMA0_Address[0] ? usedw_r : usedw_l;	
assign start_cond = (usedw >= WORDS - 1);

//Next state logic
always @ (*) begin
	NextState = CurrentState;
	case (CurrentState)
	WAIT4DMA:	begin
						if (DMA1_Ready_r && !DMA0_Address[0]) 
							NextState = DR_READ;
						else if (DMA0_Ready_r && ((start_cond) || (send_cnt > 0 && send_cnt < WORDS)) && !((send_cnt == WORDS) && WR)) 
							NextState = WRITE; 
						else if ((usedw_other >= WORDS - 1)  && (send_cnt == 0)) 
							NextState = SW_BUF;
					end	
	WRITE:		begin
						if (send_cnt >= WORDS - 1)
							if (start_cond && (usedw > usedw_other))
								NextState = WAIT4DMA;
							else
								NextState = SW_BUF;
						else if (DMA0_Watermark_r) 
							NextState = PAUSE_W;
						
					end
	PAUSE_W:		begin
						if (~DMA0_Ready_r || (lat_count == 6)) 
							NextState = WAIT4DMA;
					end
	DR_READ:		begin
						if (lat_count == 4)
							NextState = READ;
					end
	READ:			begin
						if (DMA1_Watermark_r) 
							NextState = PAUSE_R;
					end
	PAUSE_R:		begin
						if (~DMA1_Ready_r) 
							NextState = RD_CMD;
					end
	RD_CMD:		begin
						case (DATA_IN[7:0])
							GET_CFG	:	begin
												if (DMA0_Ready_r & !DMA0_Watermark_r)
													NextState = SEND_CFG;
											end
							STRT_ST	:	NextState = START_ST;
							STOP_ST	:	NextState = STP_ST;
							default	:	NextState = WAIT4DMA;
						endcase
					end
	SEND_CFG:	begin
						if (rdaddress == 'h02)
							NextState = WAIT4DMA;
					end
	START_ST:	begin
						NextState = WAIT4DMA;
					end
	STP_ST:		begin
						NextState = WAIT4DMA;
					end
	SW_BUF:		begin
						if (lat_count == 6)
							NextState = WAIT4DMA;
					end
	
	default:		NextState = WAIT4DMA;		
	endcase
end
		
//Send Cnt
always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n)
	send_cnt <= 0;
else if ((send_cnt == WORDS) || (CurrentState == SEND_CFG))
	send_cnt <= 0;
else if (CurrentState == WRITE)
	send_cnt <= send_cnt + 1'b1;

//line cnt r
always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n) 
	line_cnt_r <= 0;
else if (((send_cnt == WORDS) && (line_cnt_r == IM_Y - 1) && !DMA0_Address[0]) || !start_stream) 
	line_cnt_r <= 0;
else if ((send_cnt == WORDS) && !DMA0_Address[0]) 
	line_cnt_r <= line_cnt_r + 1'b1;
	
//line cnt l
always @ (posedge USB_CLK or negedge rst_n)
if (!rst_n) 
	line_cnt_l <= 0;
else if (((send_cnt == WORDS) && (line_cnt_l == IM_Y - 1) && DMA0_Address[0]) || !start_stream) 
	line_cnt_l <= 0;
else if ((send_cnt == WORDS) && DMA0_Address[0]) 
	line_cnt_l <= line_cnt_l + 1'b1;
	
endmodule
